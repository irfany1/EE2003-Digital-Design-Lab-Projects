module multiplication(
    input [4:0] in1,
    input [6:0] in2,
    output [11:0] out
);

assign out = in1 * in2;

endmodule